`timescale 1ns/1ps

`include "axi.vh"
`include "iob_lib.vh"
`include "iob_eth.vh"
`include "iob_eth_swreg_def.vh"

/*
 Ethernet Core
*/

module iob_eth #(
                 parameter ETH_MAC_ADDR = `ETH_MAC_ADDR
                 )
   (
    // CPU side
    input                   clk,
    input                   rst,

    input                   valid,
    output reg              ready,
    input [3:0]             wstrb,
    input [`ETH_ADDR_W-1:0] addr,
    output reg [31:0]       data_out,
    input [31:0]            data_in,

    // PHY side
    output reg              ETH_PHY_RESETN,

    // PLL
    input                   PLL_LOCKED,

    // RX
    input                   RX_CLK,
    input [3:0]             RX_DATA,
    input                   RX_DV,

    // TX
    input                   TX_CLK,
    output                  TX_EN,
    output [3:0]            TX_DATA
    );

   // registers
   // dummy
   reg [31:0]               dummy_reg;
   reg                      dummy_reg_en;
   // tx_nbytes
   reg [10:0]               tx_nbytes_reg;
   reg                      tx_nbytes_reg_en;
   // rx_nbytes
   reg [10:0]               rx_nbytes_reg;
   reg                      rx_nbytes_reg_en;
   
   // control
   reg                      send_en;
   reg                      send;

   reg                      rcv_ack_en;
   reg                      rcv_ack;

   // tx signals
   reg                      tx_wr;
   reg [1:0]                tx_ready;
   reg [1:0]                tx_clk_pll_locked;
   wire                     tx_ready_int;

   // rx signals
   reg [1:0]                rx_data_rcvd;
   wire                     rx_data_rcvd_int;
   wire[31:0]               rx_rd_data;
   reg [10:0]               rx_wr_addr_cpu[1:0];
   reg [31:0]               crc_value_cpu[1:0];
   
   // phy reset timer
   reg [19:0]               phy_rst_cnt;
   reg                      phy_clk_detected;
   reg                      phy_dv_detected;
   reg [1:0]                phy_clk_detected_sync;
   reg [1:0]                phy_dv_detected_sync;

   reg                      rst_soft_en;
   reg                      rst_soft;
   wire                     rst_int;

   // ETH CLOCK DOMAIN
   wire [8:0]               tx_rd_addr;
   wire [31:0]              tx_rd_data;

   wire [10:0]              rx_wr_addr;
   wire [7:0]               rx_wr_data;
   wire                     rx_wr;
   wire [31:0]              crc_value;

   wire [8:0]               rx_address;
   wire [8:0]               tx_address;
   wire [31:0]              tx_wr_data;
   wire                     do_tx_wr;


   assign  rx_address = addr[8:0];
   assign  tx_address = addr[8:0];
   assign  tx_wr_data = data_in;
   assign  do_tx_wr   = tx_wr;


   assign rst_int = rst_soft | rst;
   
   // SYNCHRONIZERS
   always @ (posedge clk, posedge rst_int)
     if (rst_int) begin
        tx_ready <= 0;
        tx_clk_pll_locked <= 0;
        rx_data_rcvd <= 0;
        rx_wr_addr_cpu[0] <= 0;
        rx_wr_addr_cpu[1] <= 0;
        crc_value_cpu[0] <= 0;
        crc_value_cpu[1] <= 0;
        phy_clk_detected_sync <= 0;
        phy_dv_detected_sync <= 0;
     end else begin
        tx_clk_pll_locked <= {tx_clk_pll_locked[0], PLL_LOCKED};
        tx_ready <= {tx_ready[0], tx_ready_int & ETH_PHY_RESETN & PLL_LOCKED};
        rx_data_rcvd <= {rx_data_rcvd[0], rx_data_rcvd_int & ETH_PHY_RESETN};
        rx_wr_addr_cpu[0] <= rx_wr_addr;
        rx_wr_addr_cpu[1] <= rx_wr_addr_cpu[0];
        crc_value_cpu[0] <= crc_value;
        crc_value_cpu[1] <= crc_value_cpu[0];
        phy_clk_detected_sync <= {phy_clk_detected_sync[0], phy_clk_detected};
        phy_dv_detected_sync <= {phy_dv_detected_sync[0], phy_dv_detected};
     end

   // cpu interface ready signal
   always @(posedge clk, posedge rst)
     if (rst)
       ready <= 1'b0;
     else
       ready <= valid;

   //
   // ADDRESS DECODER
   //

   // write
   always @* begin
      // defaults
      rst_soft_en = 0;
      send_en = 0;
      rcv_ack_en = 0;
      dummy_reg_en = 0;
      tx_nbytes_reg_en = 0;
      rx_nbytes_reg_en = 0;
      tx_wr = 1'b0;

      if(valid & (|wstrb))
        case (addr)
          `ETH_SEND: send_en = 1'b1;
          `ETH_RCVACK: rcv_ack_en = 1'b1;
          `ETH_DUMMY: dummy_reg_en = 1'b1;
          `ETH_TX_NBYTES: tx_nbytes_reg_en = 1'b1;
          `ETH_RX_NBYTES: rx_nbytes_reg_en = 1'b1;
          `ETH_SOFTRST: rst_soft_en  = 1'b1;
          default: tx_wr = addr[11] & 1'b1; // ETH_DATA
        endcase
   end


   // read
   always @* begin
      case (addr)
        `ETH_STATUS: data_out = {16'b0, tx_clk_pll_locked[1], rx_wr_addr_cpu[1], phy_clk_detected_sync[1], phy_dv_detected_sync[1], rx_data_rcvd[1], tx_ready[1]};
        `ETH_DUMMY: data_out = dummy_reg;
        `ETH_CRC: data_out = crc_value_cpu[1];
        `ETH_RCV_SIZE: data_out = rx_wr_addr;
        default: data_out = rx_rd_data; // ETH_DATA
      endcase
   end

   //
   // REGISTERS
   //

   // soft reset self-clearing register
   always @ (posedge clk, posedge rst)
     if (rst)
       rst_soft <= 1'b1;
     else if (rst_soft_en && !rst_soft)
       rst_soft <= 1'b1;
     else
       rst_soft <= 1'b0;

   always @ (posedge clk, posedge rst_int)
     if (rst_int) begin
        tx_nbytes_reg <= 11'd46;
        rx_nbytes_reg <= 11'd46;
        dummy_reg <= 0;
     end else if (dummy_reg_en)
       dummy_reg <= data_in;
     else if (tx_nbytes_reg_en)
       tx_nbytes_reg <= data_in[10:0];
     else if (rx_nbytes_reg_en)
       rx_nbytes_reg <= data_in[10:0];
   
   // SYNCHRONIZERS

  `IOB_F2S_SYNC(TX_CLK, send_en, send_sync, send)
  `IOB_F2S_SYNC(RX_CLK, rcv_ack_en, rck_ack_sync, rcv_ack)

   //
   // TX and RX BUFFERS
   //

   iob_ram_t2p #(
                       .DATA_W(32),
                       .ADDR_W((`ETH_ADDR_W-1)-2)
                       )
   tx_buffer
   (
    // Front-End (written by host)
      .w_clk(clk),
      .w_addr(tx_address),
      .w_en(do_tx_wr),
      .w_data(tx_wr_data),

    // Back-End (read by core)
      .r_clk(TX_CLK),
      .r_addr(tx_rd_addr),
      .r_en(1'b1),
      .r_data(tx_rd_data)
   );

   // Transform 8 bit rx data to 32 bit data to be stored in rx_buffer
   reg [8:0] stored_rx_addr;
   reg [31:0] stored_rx_data; 
   reg stored_rx_wr;

   always @(posedge RX_CLK,posedge rst)
   if(rst) begin
     stored_rx_addr <= 0;
     stored_rx_data <= 0;
     stored_rx_wr <= 1'b0;
   end else if(rx_wr) begin
     stored_rx_addr <= rx_wr_addr[10:2];
     stored_rx_data[8 * rx_wr_addr[1:0] +: 8] <= rx_wr_data;
     stored_rx_wr <= 1'b1;
   end

   iob_ram_t2p #(
                       .DATA_W(32),
                       .ADDR_W((`ETH_ADDR_W-1)-2)
                       )
   rx_buffer
   (
     // Front-End (written by core)
     .w_clk(RX_CLK),
     .w_addr(stored_rx_addr),
     .w_en(stored_rx_wr),
     .w_data(stored_rx_data),

     // Back-End (read by host)
     .r_clk(clk),
     .r_addr(rx_address),
     .r_en(1'b1),
     .r_data(rx_rd_data)
   );

   //
   // TRANSMITTER
   //

   // Transform 32 bit data from tx_buffer to 8 bit data for tx input
   reg [1:0] delayed_tx_sel;
   wire [10:0] tx_out_addr;
   
   always @(posedge TX_CLK,posedge rst_int)
     if(rst_int)
       delayed_tx_sel <= 0;
     else
       delayed_tx_sel <= tx_out_addr[1:0];

   assign tx_rd_addr = tx_out_addr[10:2];
   wire [7:0] tx_in_data = delayed_tx_sel[1] ? (delayed_tx_sel[0] ? tx_rd_data[8*3 +: 8] : tx_rd_data[8*2 +: 8]):
                                               (delayed_tx_sel[0] ? tx_rd_data[8*1 +: 8] : tx_rd_data[8*0 +: 8]);

   iob_eth_tx
     tx (
         // cpu side
         .rst     (rst_int),
         .nbytes  (tx_nbytes_reg),
         .ready   (tx_ready_int),

         // mii side
         .send    (send),
         .addr    (tx_out_addr),
         .data    (tx_in_data),
         .TX_CLK  (TX_CLK),
         .TX_EN   (TX_EN),
         .TX_DATA (TX_DATA)
         );


   //
   // RECEIVER
   //

   iob_eth_rx #(
                .ETH_MAC_ADDR(ETH_MAC_ADDR)
                )
   rx (
       // cpu side
       .rst       (rst_int),
       .data_rcvd (rx_data_rcvd_int),

       // mii side
       .rcv_ack   (rcv_ack),
       .wr        (rx_wr),
       .addr      (rx_wr_addr),
       .data      (rx_wr_data),
       .RX_CLK    (RX_CLK),
       .RX_DATA   (RX_DATA),
       .RX_DV     (RX_DV),
       .crc_value (crc_value)
       );


   //
   //  PHY RESET
   //
   
   always @ (posedge clk, posedge rst_int)
     if(rst_int) begin
        phy_rst_cnt <= 0;
        ETH_PHY_RESETN <= 0;
     end else 
`ifdef SIM // Faster for simulation
       if (phy_rst_cnt != 20'h000FF)
`else
       if (phy_rst_cnt != 20'hFFFFF)
`endif
         phy_rst_cnt <= phy_rst_cnt+1'b1;
       else
         ETH_PHY_RESETN <= 1;

   reg [1:0] rx_rst;
   always @ (posedge RX_CLK, negedge ETH_PHY_RESETN)
     if (!ETH_PHY_RESETN)
       rx_rst <= 2'b11;
     else
       rx_rst <= {rx_rst[0], 1'b0};
   
   always @ (posedge RX_CLK, posedge rx_rst[1])
     if (rx_rst[1]) begin
        phy_clk_detected <= 1'b0;
        phy_dv_detected <= 1'b0;
     end else begin 
        phy_clk_detected <= 1'b1;
        if(RX_DV)
          phy_dv_detected <= 1'b1;
     end

endmodule
