`define SFD 8'hD5
`define MAC_ADDR 48'h00aa0062c606
