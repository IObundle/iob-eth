// The SWREGs are defined manually in iob_eth.v
// this file exists for correct integration in iob-soc type systems
