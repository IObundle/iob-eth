// SPDX-FileCopyrightText: 2025 IObundle
//
// SPDX-License-Identifier: MIT

`include "iob_eth_csrs_conf.vh"
`define IOB_CSRS_ADDR_W (`IOB_ETH_CSRS_ADDR_W+2)
