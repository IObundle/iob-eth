// SPDX-FileCopyrightText: 2025 IObundle
//
// SPDX-License-Identifier: MIT

// megafunction wizard: %altddio_out%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTDDIO_OUT 

// ============================================================
// File Name: ddio_out_clkbuf.v
// Megafunction Name(s):
// 			ALTDDIO_OUT
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 20.1.0 Build 711 06/05/2020 SJ Standard Edition
// ************************************************************



// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module ddio_out_clkbuf (
   aclr,
   datain_h,
   datain_l,
   outclock,
   dataout
);

   input aclr;
   input [0:0] datain_h;
   input [0:0] datain_l;
   input outclock;
   output [0:0] dataout;

   wire [0:0] sub_wire0;
   wire [0:0] dataout = sub_wire0[0:0];

   altddio_out ALTDDIO_OUT_component (
      .aclr      (aclr),
      .datain_h  (datain_h),
      .datain_l  (datain_l),
      .outclock  (outclock),
      .dataout   (sub_wire0),
      .aset      (1'b0),
      .oe        (1'b1),
      .oe_out    (),
      .outclocken(1'b1),
      .sclr      (1'b0),
      .sset      (1'b0)
   );
   defparam ALTDDIO_OUT_component.extend_oe_disable = "OFF",
       ALTDDIO_OUT_component.intended_device_family = "Cyclone V",
       ALTDDIO_OUT_component.invert_output = "OFF", ALTDDIO_OUT_component.lpm_hint = "UNUSED",
       ALTDDIO_OUT_component.lpm_type = "altddio_out", ALTDDIO_OUT_component.oe_reg =
       "UNREGISTERED", ALTDDIO_OUT_component.power_up_high = "OFF", ALTDDIO_OUT_component.width = 1;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: EXTEND_OE_DISABLE STRING "OFF"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: INVERT_OUTPUT STRING "OFF"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altddio_out"
// Retrieval info: CONSTANT: OE_REG STRING "UNREGISTERED"
// Retrieval info: CONSTANT: POWER_UP_HIGH STRING "OFF"
// Retrieval info: CONSTANT: WIDTH NUMERIC "1"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: USED_PORT: datain_h 0 0 1 0 INPUT NODEFVAL "datain_h[0..0]"
// Retrieval info: CONNECT: @datain_h 0 0 1 0 datain_h 0 0 1 0
// Retrieval info: USED_PORT: datain_l 0 0 1 0 INPUT NODEFVAL "datain_l[0..0]"
// Retrieval info: CONNECT: @datain_l 0 0 1 0 datain_l 0 0 1 0
// Retrieval info: USED_PORT: dataout 0 0 1 0 OUTPUT NODEFVAL "dataout[0..0]"
// Retrieval info: CONNECT: dataout 0 0 1 0 @dataout 0 0 1 0
// Retrieval info: USED_PORT: outclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL "outclock"
// Retrieval info: CONNECT: @outclock 0 0 0 0 outclock 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL ddio_out_clkbuf.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ddio_out_clkbuf.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ddio_out_clkbuf.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ddio_out_clkbuf_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ddio_out_clkbuf_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ddio_out_clkbuf.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ddio_out_clkbuf.cmp TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ddio_out_clkbuf.ppf TRUE FALSE
// Retrieval info: LIB_FILE: altera_mf
