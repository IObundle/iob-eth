    // TX Front-End
    .iob_eth_tx_buffer_enA(iob_eth_tx_buffer_enA),
    .iob_eth_tx_buffer_weA(iob_eth_tx_buffer_weA),
    .iob_eth_tx_buffer_addrA(iob_eth_tx_buffer_addrA),
    .iob_eth_tx_buffer_dinA(iob_eth_tx_buffer_dinA),
    // TX Back-End
    .iob_eth_tx_buffer_addrB(iob_eth_tx_buffer_addrB),
    .iob_eth_tx_buffer_doutB(iob_eth_tx_buffer_doutB),
    // RX Front-End
    .iob_eth_rx_buffer_enA(iob_eth_rx_buffer_enA),
    .iob_eth_rx_buffer_weA(iob_eth_rx_buffer_weA),
    .iob_eth_rx_buffer_addrA(iob_eth_rx_buffer_addrA),
    .iob_eth_rx_buffer_dinA(iob_eth_rx_buffer_dinA),
    // RX Back-End
    .iob_eth_rx_buffer_enB(iob_eth_rx_buffer_enB),
    .iob_eth_rx_buffer_addrB(iob_eth_rx_buffer_addrB),
    .iob_eth_rx_buffer_doutB(iob_eth_rx_buffer_doutB),
